`timescale 1ns / 1ns

module tb_bram();

   reg clk_l;
   reg rst_n;

   parameter CLK_PERIOD = 200;
   parameter WID_W = 16;
   parameter WID_WADDR = 10;   

   initial begin
      clk_l = 1'b1;
      forever #(CLK_PERIOD/2) clk_l = ~clk_l;
   end

   initial begin
      rst_n = 1'b1;
      repeat(2) @(negedge clk_l);
      rst_n = 1'b0;
      repeat(20) @(negedge clk_l);
      rst_n = 1'b1;
   end

   reg [WID_WADDR-1:0] w_rd_addr;
   wire [WID_W-1:0] w_rd_data;

   initial begin
      forever begin
         @(posedge clk_l);
         if(~rst_n) begin
            w_rd_addr <= 0;
         end else begin
            w_rd_addr <= w_rd_addr + 1;
         end
      end
   end
 
   RAMB18E2 #(
      // CASCADE_ORDER_A, CASCADE_ORDER_B: "FIRST", "MIDDLE", "LAST", "NONE" 
      .CASCADE_ORDER_A("NONE"),
      .CASCADE_ORDER_B("NONE"),
      // CLOCK_DOMAINS: "COMMON", "INDEPENDENT" 
      .CLOCK_DOMAINS("INDEPENDENT"),
      // Collision check: "ALL", "GENERATE_X_ONLY", "NONE", "WARNING_ONLY" 
      .SIM_COLLISION_CHECK("ALL"),
      // DOA_REG, DOB_REG: Optional output register (0, 1)
      .DOA_REG(1),
      // .DOB_REG(1),
      // ENADDRENA/ENADDRENB: Address enable pin enable, "TRUE", "FALSE" 
      .ENADDRENA("FALSE"),
      .ENADDRENB("FALSE"),
      // INITP_00 to INITP_07: Initial contents of parity memory array
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // INIT_00 to INIT_3F: Initial contents of data memory array
      .INIT_00(256'hdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddd),
      .INIT_01(256'hdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddd),
      .INIT_02(256'hdddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddd),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // INIT_A, INIT_B: Initial values on output ports
      .INIT_A(18'h00000),
      .INIT_B(18'h00000),
      // Initialization File: RAM initialization file
      .INIT_FILE("NONE"),
      // Programmable Inversion Attributes: Specifies the use of the built-in programmable inversion
      .IS_CLKARDCLK_INVERTED(1'b0),
      .IS_CLKBWRCLK_INVERTED(1'b0),
      .IS_ENARDEN_INVERTED(1'b0),
      .IS_ENBWREN_INVERTED(1'b0),
      .IS_RSTRAMARSTRAM_INVERTED(1'b0),
      .IS_RSTRAMB_INVERTED(1'b0),
      .IS_RSTREGARSTREG_INVERTED(1'b0),
      .IS_RSTREGB_INVERTED(1'b0),
      // RDADDRCHANGE: Disable memory access when output value does not change ("TRUE", "FALSE")
      .RDADDRCHANGEA("FALSE"),
      .RDADDRCHANGEB("FALSE"),
      // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
      .READ_WIDTH_A(18),                                                                 // 0-9
      .READ_WIDTH_B(0),                                                                 // 0-9
      .WRITE_WIDTH_A(0),                                                                // 0-9
      .WRITE_WIDTH_B(0),                                                                // 0-9
      // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG", "REGCE")
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      // SRVAL_A, SRVAL_B: Set/reset value for output
      .SRVAL_A(18'h00000),
      .SRVAL_B(18'h00000),
      // Sleep Async: Sleep function asynchronous or synchronous ("TRUE", "FALSE")
      .SLEEP_ASYNC("FALSE"),
      // WriteMode: "WRITE_FIRST", "NO_CHANGE", "READ_FIRST" 
      .WRITE_MODE_A("READ_FIRST"),
      .WRITE_MODE_B("READ_FIRST") 
   )
   RAMB18E2_inst (
      // Cascade Signals outputs: Multi-BRAM cascade signals
      // .CASDOUTA(CASDOUTA),               // 16-bit output: Port A cascade output data
      // .CASDOUTB(CASDOUTB),               // 16-bit output: Port B cascade output data
      // .CASDOUTPA(CASDOUTPA),             // 2-bit output: Port A cascade output parity data
      // .CASDOUTPB(CASDOUTPB),             // 2-bit output: Port B cascade output parity data
      // Port A Data outputs: Port A data
      .DOUTADOUT(w_rd_data),             // 16-bit output: Port A data/LSB data
      // .DOUTPADOUTP(DOUTPADOUTP),         // 2-bit output: Port A parity/LSB parity
      // Port B Data outputs: Port B data
      // .DOUTBDOUT(DOUTBDOUT),             // 16-bit output: Port B data/MSB data
      // .DOUTPBDOUTP(DOUTPBDOUTP),         // 2-bit output: Port B parity/MSB parity
      // Cascade Signals inputs: Multi-BRAM cascade signals
      // .CASDIMUXA(CASDIMUXA),             // 1-bit input: Port A input data (0=DINA, 1=CASDINA)
      // .CASDIMUXB(CASDIMUXB),             // 1-bit input: Port B input data (0=DINB, 1=CASDINB)
      // .CASDINA(CASDINA),                 // 16-bit input: Port A cascade input data
      // .CASDINB(CASDINB),                 // 16-bit input: Port B cascade input data
      // .CASDINPA(CASDINPA),               // 2-bit input: Port A cascade input parity data
      // .CASDINPB(CASDINPB),               // 2-bit input: Port B cascade input parity data
      // .CASDOMUXA(CASDOMUXA),             // 1-bit input: Port A unregistered data (0=BRAM data, 1=CASDINA)
      // .CASDOMUXB(CASDOMUXB),             // 1-bit input: Port B unregistered data (0=BRAM data, 1=CASDINB)
      // .CASDOMUXEN_A(CASDOMUXEN_A),       // 1-bit input: Port A unregistered output data enable
      // .CASDOMUXEN_B(CASDOMUXEN_B),       // 1-bit input: Port B unregistered output data enable
      // .CASOREGIMUXA(CASOREGIMUXA),       // 1-bit input: Port A registered data (0=BRAM data, 1=CASDINA)
      // .CASOREGIMUXB(CASOREGIMUXB),       // 1-bit input: Port B registered data (0=BRAM data, 1=CASDINB)
      // .CASOREGIMUXEN_A(CASOREGIMUXEN_A), // 1-bit input: Port A registered output data enable
      // .CASOREGIMUXEN_B(CASOREGIMUXEN_B), // 1-bit input: Port B registered output data enable
      // Port A Address/Control Signals inputs: Port A address and control signals
      .ADDRARDADDR({w_rd_addr, 4'b0000}),         // 14-bit input: A/Read port address
      .ADDRENA(1'b1),                 // 1-bit input: Active-High A/Read port address enable
      .CLKARDCLK(clk_l),             // 1-bit input: A/Read port clock
      .ENARDEN(1'b1),                 // 1-bit input: Port A enable/Read enable
      .REGCEAREGCE(1'b1),         // 1-bit input: Port A register enable/Register enable
      .RSTRAMARSTRAM(~rst_n),     // 1-bit input: Port A set/reset
      .RSTREGARSTREG(~rst_n),     // 1-bit input: Port A register set/reset
      .WEA(2'b00)                         // 2-bit input: Port A write enable
      // Port A Data inputs: Port A data
      // .DINADIN(DINADIN),                 // 16-bit input: Port A data/LSB data
      // .DINPADINP(DINPADINP),             // 2-bit input: Port A parity/LSB parity
      // Port B Address/Control Signals inputs: Port B address and control signals
      // .ADDRBWRADDR(ADDRBWRADDR),         // 14-bit input: B/Write port address
      // .ADDRENB(ADDRENB),                 // 1-bit input: Active-High B/Write port address enable
      // .CLKBWRCLK(CLKBWRCLK),             // 1-bit input: B/Write port clock
      // .ENBWREN(ENBWREN),                 // 1-bit input: Port B enable/Write enable
      // .REGCEB(REGCEB),                   // 1-bit input: Port B register enable
      // .RSTRAMB(RSTRAMB),                 // 1-bit input: Port B set/reset
      // .RSTREGB(RSTREGB),                 // 1-bit input: Port B register set/reset
      // .SLEEP(SLEEP),                     // 1-bit input: Sleep Mode
      // .WEBWE(WEBWE),                     // 4-bit input: Port B write enable/Write enable
      // Port B Data inputs: Port B data
      // .DINBDIN(DINBDIN),                 // 16-bit input: Port B data/MSB data
      // .DINPBDINP(DINPBDINP)              // 2-bit input: Port B parity/MSB parity
   );





endmodule // tb_bram










